library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MaqEstados_testbench2 is
end MaqEstados_testbench2;

architecture MaqEstados_TB_arch of MaqEstados_testbench2 is

-- Component Declaration
component Maq_estados
    port (
        clk, front_sensor, back_sensor, cobrar, reset: in std_logic;
        cat: in std_logic_vector(1 downto 0);
        id: in std_logic_vector(2 downto 0);
        tala_ini, tala_fin, alar_son, led, sema_ini, sema_fin, cont_vehiculo: out std_logic;
        contador: buffer integer range 0 to 2
    );
end component;

-- Signals Declaration
signal clk_TB, front_sensor_TB, back_sensor_TB, cobrar_TB, reset_TB: std_logic := '0';
signal cat_TB: std_logic_vector(1 downto 0) := "00";
signal id_TB: std_logic_vector(2 downto 0) := "000";
signal tala_ini_TB, tala_fin_TB, alar_son_TB, led_TB, sema_ini_TB, sema_fin_TB, cont_vehiculo_TB: std_logic;
signal contador_TB: integer := 0;

begin

-- DUT Instantiation
DUT1: Maq_estados
    port map (
        clk => clk_TB,
        front_sensor => front_sensor_TB,
        back_sensor => back_sensor_TB,
        cobrar => cobrar_TB,
        reset => reset_TB,
        cat => cat_TB,
        id => id_TB,
        tala_ini => tala_ini_TB,
        tala_fin => tala_fin_TB,
        alar_son => alar_son_TB,
        led => led_TB,
        sema_ini => sema_ini_TB,
        sema_fin => sema_fin_TB,
        cont_vehiculo => cont_vehiculo_TB,
        contador => contador_TB
    );

-- Stimulus Generation
STIMULUS: process
begin
    -- Reset inicial
    reset_TB <= '1';
    wait for 10 ns;
    reset_TB <= '0';
    wait for 10 ns;

    -- Prueba del estado "Inicio"
    front_sensor_TB <= '1';
    back_sensor_TB <= '1';
    cat_TB <= "01";
    id_TB <= "001";
    wait for 10 ns;

    -- Prueba del estado "Identificador de vehículo"
    cat_TB <= "00"; -- Rojo
    wait for 10 ns;
    cat_TB <= "01"; -- Verde
    wait for 10 ns;

    -- Prueba del estado "Incorrecta"
    id_TB <= "000";
    wait for 10 ns;
    id_TB <= "010";
    wait for 10 ns;

    -- Prueba del estado "Realizar Cobro"
    id_TB <= "001";
    cobrar_TB <= '1';
    wait for 10 ns;
    cobrar_TB <= '0';
    wait for 10 ns;

    -- Prueba de salida "Salida"
    wait for 10 ns;

    -- Reinicio de la máquina de estados
    reset_TB <= '1';
    wait for 10 ns;
    reset_TB <= '0';
    wait for 10 ns;

    -- Caso 1: Probar la transición al estado "Incorrecta" cuando el identificador es inválido y la categoría es roja
    cat_TB <= "00"; -- Rojo
    id_TB <= "101"; -- Identificador inválido
    wait for 10 ns;

    -- Caso 2: Probar la transición desde "Realizar Cobro" a "Salida" cuando se realiza el cobro correctamente
    id_TB <= "001"; -- Identificador válido
    cobrar_TB <= '1';
    wait for 10 ns;
    cobrar_TB <= '0';
    wait for 20 ns; -- Tiempo adicional para permitir la transición a "Salida"

    -- Caso 3: Probar la transición desde "Inicio" a "Identificador de vehículo" cuando la categoría es roja
    front_sensor_TB <= '1';
    back_sensor_TB <= '1';
    cat_TB <= "00"; -- Rojo
    id_TB <= "001"; -- Identificador válido
    wait for 10 ns;

    -- Caso 4: Probar la transición desde "Identificador de vehículo" a "Incorrecta" cuando el identificador es inválido y la categoría es verde
    cat_TB <= "01"; -- Verde
    id_TB <= "111"; -- Identificador inválido
    wait for 10 ns;

    -- Caso 5: Probar la transición desde "Realizar Cobro" a "Inicio" después de realizar el cobro correctamente
    id_TB <= "001"; -- Identificador válido
    cobrar_TB <= '1';
    wait for 10 ns;
    cobrar_TB <= '0';
    wait for 20 ns; -- Tiempo adicional para permitir la transición a "Salida"
    front_sensor_TB <= '1';
    back_sensor_TB <= '1';
    cat_TB <= "01"; -- Verde
    id_TB <= "001"; -- Identificador válido
    wait for 10 ns;

    wait; -- Espera indefinidamente
end process STIMULUS;

end MaqEstados_TB_arch;